magic
tech sky130A
magscale 1 2
timestamp 1710672453
<< obsli1 >>
rect 1104 2159 38824 597329
<< obsm1 >>
rect 934 2128 38824 597360
<< metal2 >>
rect 9954 0 10010 800
rect 29918 0 29974 800
<< obsm2 >>
rect 938 856 35242 597349
rect 938 800 9898 856
rect 10066 800 29862 856
rect 30030 800 35242 856
<< metal3 >>
rect 0 586984 800 587104
rect 0 569032 800 569152
rect 0 551080 800 551200
rect 0 533128 800 533248
rect 0 515176 800 515296
rect 0 497224 800 497344
rect 0 479272 800 479392
rect 0 461320 800 461440
rect 0 443368 800 443488
rect 0 425416 800 425536
rect 0 407464 800 407584
rect 0 389512 800 389632
rect 0 371560 800 371680
rect 0 353608 800 353728
rect 0 335656 800 335776
rect 0 317704 800 317824
rect 0 299752 800 299872
rect 0 281800 800 281920
rect 0 263848 800 263968
rect 0 245896 800 246016
rect 0 227944 800 228064
rect 0 209992 800 210112
rect 0 192040 800 192160
rect 0 174088 800 174208
rect 0 156136 800 156256
rect 0 138184 800 138304
rect 0 120232 800 120352
rect 0 102280 800 102400
rect 0 84328 800 84448
rect 0 66376 800 66496
rect 0 48424 800 48544
rect 0 30472 800 30592
rect 0 12520 800 12640
<< obsm3 >>
rect 800 587184 35246 597345
rect 880 586904 35246 587184
rect 800 569232 35246 586904
rect 880 568952 35246 569232
rect 800 551280 35246 568952
rect 880 551000 35246 551280
rect 800 533328 35246 551000
rect 880 533048 35246 533328
rect 800 515376 35246 533048
rect 880 515096 35246 515376
rect 800 497424 35246 515096
rect 880 497144 35246 497424
rect 800 479472 35246 497144
rect 880 479192 35246 479472
rect 800 461520 35246 479192
rect 880 461240 35246 461520
rect 800 443568 35246 461240
rect 880 443288 35246 443568
rect 800 425616 35246 443288
rect 880 425336 35246 425616
rect 800 407664 35246 425336
rect 880 407384 35246 407664
rect 800 389712 35246 407384
rect 880 389432 35246 389712
rect 800 371760 35246 389432
rect 880 371480 35246 371760
rect 800 353808 35246 371480
rect 880 353528 35246 353808
rect 800 335856 35246 353528
rect 880 335576 35246 335856
rect 800 317904 35246 335576
rect 880 317624 35246 317904
rect 800 299952 35246 317624
rect 880 299672 35246 299952
rect 800 282000 35246 299672
rect 880 281720 35246 282000
rect 800 264048 35246 281720
rect 880 263768 35246 264048
rect 800 246096 35246 263768
rect 880 245816 35246 246096
rect 800 228144 35246 245816
rect 880 227864 35246 228144
rect 800 210192 35246 227864
rect 880 209912 35246 210192
rect 800 192240 35246 209912
rect 880 191960 35246 192240
rect 800 174288 35246 191960
rect 880 174008 35246 174288
rect 800 156336 35246 174008
rect 880 156056 35246 156336
rect 800 138384 35246 156056
rect 880 138104 35246 138384
rect 800 120432 35246 138104
rect 880 120152 35246 120432
rect 800 102480 35246 120152
rect 880 102200 35246 102480
rect 800 84528 35246 102200
rect 880 84248 35246 84528
rect 800 66576 35246 84248
rect 880 66296 35246 66576
rect 800 48624 35246 66296
rect 880 48344 35246 48624
rect 800 30672 35246 48344
rect 880 30392 35246 30672
rect 800 12720 35246 30392
rect 880 12440 35246 12720
rect 800 2143 35246 12440
<< metal4 >>
rect 4208 2128 4528 597360
rect 19568 2128 19888 597360
rect 34928 2128 35248 597360
<< obsm4 >>
rect 1531 167043 4128 353429
rect 4608 167043 7669 353429
<< labels >>
rlabel metal3 s 0 586984 800 587104 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 48424 800 48544 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 533128 800 533248 6 io_in[1]
port 3 nsew signal input
rlabel metal3 s 0 479272 800 479392 6 io_in[2]
port 4 nsew signal input
rlabel metal3 s 0 425416 800 425536 6 io_in[3]
port 5 nsew signal input
rlabel metal3 s 0 371560 800 371680 6 io_in[4]
port 6 nsew signal input
rlabel metal3 s 0 317704 800 317824 6 io_in[5]
port 7 nsew signal input
rlabel metal3 s 0 263848 800 263968 6 io_in[6]
port 8 nsew signal input
rlabel metal3 s 0 209992 800 210112 6 io_in[7]
port 9 nsew signal input
rlabel metal3 s 0 156136 800 156256 6 io_in[8]
port 10 nsew signal input
rlabel metal3 s 0 102280 800 102400 6 io_in[9]
port 11 nsew signal input
rlabel metal3 s 0 551080 800 551200 6 io_oeb[0]
port 12 nsew signal output
rlabel metal3 s 0 12520 800 12640 6 io_oeb[10]
port 13 nsew signal output
rlabel metal3 s 0 497224 800 497344 6 io_oeb[1]
port 14 nsew signal output
rlabel metal3 s 0 443368 800 443488 6 io_oeb[2]
port 15 nsew signal output
rlabel metal3 s 0 389512 800 389632 6 io_oeb[3]
port 16 nsew signal output
rlabel metal3 s 0 335656 800 335776 6 io_oeb[4]
port 17 nsew signal output
rlabel metal3 s 0 281800 800 281920 6 io_oeb[5]
port 18 nsew signal output
rlabel metal3 s 0 227944 800 228064 6 io_oeb[6]
port 19 nsew signal output
rlabel metal3 s 0 174088 800 174208 6 io_oeb[7]
port 20 nsew signal output
rlabel metal3 s 0 120232 800 120352 6 io_oeb[8]
port 21 nsew signal output
rlabel metal3 s 0 66376 800 66496 6 io_oeb[9]
port 22 nsew signal output
rlabel metal3 s 0 569032 800 569152 6 io_out[0]
port 23 nsew signal output
rlabel metal3 s 0 30472 800 30592 6 io_out[10]
port 24 nsew signal output
rlabel metal3 s 0 515176 800 515296 6 io_out[1]
port 25 nsew signal output
rlabel metal3 s 0 461320 800 461440 6 io_out[2]
port 26 nsew signal output
rlabel metal3 s 0 407464 800 407584 6 io_out[3]
port 27 nsew signal output
rlabel metal3 s 0 353608 800 353728 6 io_out[4]
port 28 nsew signal output
rlabel metal3 s 0 299752 800 299872 6 io_out[5]
port 29 nsew signal output
rlabel metal3 s 0 245896 800 246016 6 io_out[6]
port 30 nsew signal output
rlabel metal3 s 0 192040 800 192160 6 io_out[7]
port 31 nsew signal output
rlabel metal3 s 0 138184 800 138304 6 io_out[8]
port 32 nsew signal output
rlabel metal3 s 0 84328 800 84448 6 io_out[9]
port 33 nsew signal output
rlabel metal4 s 4208 2128 4528 597360 6 vccd1
port 34 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 597360 6 vccd1
port 34 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 597360 6 vssd1
port 35 nsew ground bidirectional
rlabel metal2 s 9954 0 10010 800 6 wb_clk_i
port 36 nsew signal input
rlabel metal2 s 29918 0 29974 800 6 wb_rst_i
port 37 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 40000 600000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7799620
string GDS_FILE /home/nihar/rvcorep_caravel/openlane/user_proj_timer/runs/24_03_17_16_13/results/signoff/user_proj_timer.magic.gds
string GDS_START 413042
<< end >>

